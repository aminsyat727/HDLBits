module top_module( output one );

// Insert your code here
    assign one = 32'h00000001;

endmodule
